
 downto 0

std_logic