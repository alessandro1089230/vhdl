
 downto 0

std_logic
15 downto 0